library verilog;
use verilog.vl_types.all;
entity register_file_vlg_vec_tst is
end register_file_vlg_vec_tst;
